[build-menu]
FT_01_LB=Compile
FT_01_CM=ghdl -a "%f" && ghdl -e "%e"
FT_01_WD=
EX_00_LB=_Execute
EX_00_CM="./%e"
EX_00_WD=
